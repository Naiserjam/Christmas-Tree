// Copyright (C) 1991-2009 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// Generated by Quartus II Version 9.1 Build 222 10/21/2009 SJ Web Edition
// Created on Tue Dec 12 17:08:24 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module final1 (
    reset,clock,dir,
    AA20,AB20,AB19,AA18,AB17,W17,T15,V15,AB9,AA9,AB7,R14,T9,R12,T10);

    input reset;
    input clock;
    input dir;
    tri0 reset;
    tri0 dir;
    output AA20;
    output AB20;
    output AB19;
    output AA18;
    output AB17;
    output W17;
    output T15;
    output V15;
    output AB9;
    output AA9;
    output AB7;
    output R14;
    output T9;
    output R12;
    output T10;
    reg AA20;
    reg reg_AA20;
    reg AB20;
    reg reg_AB20;
    reg AB19;
    reg reg_AB19;
    reg AA18;
    reg reg_AA18;
    reg AB17;
    reg reg_AB17;
    reg W17;
    reg reg_W17;
    reg T15;
    reg reg_T15;
    reg V15;
    reg reg_V15;
    reg AB9;
    reg reg_AB9;
    reg AA9;
    reg reg_AA9;
    reg AB7;
    reg reg_AB7;
    reg R14;
    reg reg_R14;
    reg T9;
    reg reg_T9;
    reg R12;
    reg reg_R12;
    reg T10;
    reg reg_T10;
    reg [14:0] fstate;
    reg [14:0] reg_fstate;
    parameter state1=0,state2=1,state3=2,state4=3,state5=4,state6=5,state7=6,state8=7,state9=8,state10=9,state11=10,state12=11,state13=12,state14=13,state15=14;

    initial
    begin
        reg_AA20 <= 1'b0;
        reg_AB20 <= 1'b0;
        reg_AB19 <= 1'b0;
        reg_AA18 <= 1'b0;
        reg_AB17 <= 1'b0;
        reg_W17 <= 1'b0;
        reg_T15 <= 1'b0;
        reg_V15 <= 1'b0;
        reg_AB9 <= 1'b0;
        reg_AA9 <= 1'b0;
        reg_AB7 <= 1'b0;
        reg_R14 <= 1'b0;
        reg_T9 <= 1'b0;
        reg_R12 <= 1'b0;
        reg_T10 <= 1'b0;
    end

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
            AA20 <= reg_AA20;
            AB20 <= reg_AB20;
            AB19 <= reg_AB19;
            AA18 <= reg_AA18;
            AB17 <= reg_AB17;
            W17 <= reg_W17;
            T15 <= reg_T15;
            V15 <= reg_V15;
            AB9 <= reg_AB9;
            AA9 <= reg_AA9;
            AB7 <= reg_AB7;
            R14 <= reg_R14;
            T9 <= reg_T9;
            R12 <= reg_R12;
            T10 <= reg_T10;
        end
    end

    always @(fstate or reset or dir)
    begin
        if (~reset) begin
            reg_fstate <= state1;
            reg_AA20 <= 1'b0;
            reg_AB20 <= 1'b0;
            reg_AB19 <= 1'b0;
            reg_AA18 <= 1'b0;
            reg_AB17 <= 1'b0;
            reg_W17 <= 1'b0;
            reg_T15 <= 1'b0;
            reg_V15 <= 1'b0;
            reg_AB9 <= 1'b0;
            reg_AA9 <= 1'b0;
            reg_AB7 <= 1'b0;
            reg_R14 <= 1'b0;
            reg_T9 <= 1'b0;
            reg_R12 <= 1'b0;
            reg_T10 <= 1'b0;
        end
        else begin
            reg_AA20 <= 1'b0;
            reg_AB20 <= 1'b0;
            reg_AB19 <= 1'b0;
            reg_AA18 <= 1'b0;
            reg_AB17 <= 1'b0;
            reg_W17 <= 1'b0;
            reg_T15 <= 1'b0;
            reg_V15 <= 1'b0;
            reg_AB9 <= 1'b0;
            reg_AA9 <= 1'b0;
            reg_AB7 <= 1'b0;
            reg_R14 <= 1'b0;
            reg_T9 <= 1'b0;
            reg_R12 <= 1'b0;
            reg_T10 <= 1'b0;
            case (fstate)
                state1: begin
                    if (dir)
                        reg_fstate <= state2;
                    else if (~(dir))
                        reg_fstate <= state15;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    reg_AA20 <= 1'b1;
                end
                state2: begin
                    if (dir)
                        reg_fstate <= state3;
                    else if (~(dir))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    reg_W17 <= 1'b1;

                    reg_AB20 <= 1'b1;
                end
                state3: begin
                    if (dir)
                        reg_fstate <= state4;
                    else if (~(dir))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    reg_AB19 <= 1'b1;

                    reg_T15 <= 1'b1;

                    reg_AA9 <= 1'b1;
                end
                state4: begin
                    if (dir)
                        reg_fstate <= state5;
                    else if (~(dir))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state4;

                    reg_AA18 <= 1'b1;

                    reg_AB7 <= 1'b1;

                    reg_V15 <= 1'b1;

                    reg_T9 <= 1'b1;
                end
                state5: begin
                    if (dir)
                        reg_fstate <= state6;
                    else if (~(dir))
                        reg_fstate <= state4;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state5;

                    reg_AB17 <= 1'b1;

                    reg_AB9 <= 1'b1;

                    reg_R14 <= 1'b1;

                    reg_T10 <= 1'b1;

                    reg_R12 <= 1'b1;
                end
                state6: begin
                    if (dir)
                        reg_fstate <= state7;
                    else if (~(dir))
                        reg_fstate <= state5;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state6;

                    reg_AB17 <= 1'b1;
                end
                state7: begin
                    if (dir)
                        reg_fstate <= state8;
                    else if (~(dir))
                        reg_fstate <= state6;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state7;

                    reg_AB9 <= 1'b1;

                    reg_AA18 <= 1'b1;
                end
                state8: begin
                    if (dir)
                        reg_fstate <= state9;
                    else if (~(dir))
                        reg_fstate <= state7;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state8;

                    reg_R14 <= 1'b1;

                    reg_V15 <= 1'b1;

                    reg_AB19 <= 1'b1;
                end
                state9: begin
                    if (dir)
                        reg_fstate <= state10;
                    else if (~(dir))
                        reg_fstate <= state8;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state9;

                    reg_AB7 <= 1'b1;

                    reg_R12 <= 1'b1;

                    reg_T15 <= 1'b1;

                    reg_AB20 <= 1'b1;
                end
                state10: begin
                    if (dir)
                        reg_fstate <= state11;
                    else if (~(dir))
                        reg_fstate <= state9;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state10;

                    reg_T10 <= 1'b1;

                    reg_W17 <= 1'b1;

                    reg_AA9 <= 1'b1;

                    reg_T9 <= 1'b1;

                    reg_AA20 <= 1'b1;
                end
                state11: begin
                    if (dir)
                        reg_fstate <= state12;
                    else if (~(dir))
                        reg_fstate <= state10;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state11;

                    reg_AB17 <= 1'b1;

                    reg_AA18 <= 1'b1;

                    reg_AB19 <= 1'b1;

                    reg_AA20 <= 1'b1;

                    reg_AB20 <= 1'b1;
                end
                state12: begin
                    if (dir)
                        reg_fstate <= state13;
                    else if (~(dir))
                        reg_fstate <= state11;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state12;

                    reg_AB9 <= 1'b1;

                    reg_V15 <= 1'b1;

                    reg_W17 <= 1'b1;

                    reg_T15 <= 1'b1;
                end
                state13: begin
                    if (dir)
                        reg_fstate <= state14;
                    else if (~(dir))
                        reg_fstate <= state12;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state13;

                    reg_R14 <= 1'b1;

                    reg_AB7 <= 1'b1;

                    reg_AA9 <= 1'b1;
                end
                state14: begin
                    if (dir)
                        reg_fstate <= state15;
                    else if (~(dir))
                        reg_fstate <= state13;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state14;

                    reg_R12 <= 1'b1;

                    reg_T9 <= 1'b1;
                end
                state15: begin
                    if (dir)
                        reg_fstate <= state1;
                    else if (~(dir))
                        reg_fstate <= state14;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state15;

                    reg_T10 <= 1'b1;
                end
                default: begin
                    reg_AA20 <= 1'bx;
                    reg_AB20 <= 1'bx;
                    reg_AB19 <= 1'bx;
                    reg_AA18 <= 1'bx;
                    reg_AB17 <= 1'bx;
                    reg_W17 <= 1'bx;
                    reg_T15 <= 1'bx;
                    reg_V15 <= 1'bx;
                    reg_AB9 <= 1'bx;
                    reg_AA9 <= 1'bx;
                    reg_AB7 <= 1'bx;
                    reg_R14 <= 1'bx;
                    reg_T9 <= 1'bx;
                    reg_R12 <= 1'bx;
                    reg_T10 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // final1
